`timescale 1 ns / 100 ps

module FourModeTimer_tb;
	reg clk;
	reg set_n;
	reg hold;
	reg C1;
	reg C2;
	
	wire [6:0] Hex_M1;
	wire [6:0] Hex_M2;
	wire [6:0] Hex_S1;
	wire [6:0] Hex_S2;
	wire CLK_ind;
	
	
endmodule
