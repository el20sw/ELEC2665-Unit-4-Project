`timescale 1 ns / 100 ps

module TimerLogic_tb;	//testbench for the the timer logic module
	reg clk_1Hz;
	reg set_n;
	reg hold;
	reg [5:0] Qs_set;
	reg [1:0] Qm_set;

	wire [5:0] Qs;
	wire [1:0] Qm;

	
	
endmodule
