`timescale 1 ns / 100 ps

module SevenSegEncoder_tb;		//testbench for the the SevenSegEncoder module
	
	reg [5:0] Qs;
	reg [1:0] Qm;
	
	wire [6:0] HexM_1;
	wire [6:0] HexM_2;
	wire [6:0] HexS_1;
	wire [6:0] HexS_2;

	
	
endmodule
